`ifndef GUARD_REGMODEL
`define GUARD_REGMODEL

bit [7:0] length_reg_copy = 0;
bit [7:0] max_burst_size_reg_copy= 0;

int errors = 0;

`endif
